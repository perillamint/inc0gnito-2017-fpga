// Reading file 'inc0gnito.asc'..

module chip (output \data[18] , output \data[17] , output \data[14] , output \data[11] , output \data[10] , output \data[6] , output \data[2] , output \data[0] , output \data[22] , output \data[16] , output \data[15] , output \data[13] , output \data[12] , output \data[9] , output \data[8] , output \data[7] , output \data[5] , output \data[4] , output \data[3] , output \data[1] , input \key[31] , input \key[30] , input \key[29] , input \key[28] , input \key[27] , input \key[26] , input \key[25] , input \key[24] , input \key[23] , input \key[22] , input \key[21] , input \key[20] , input \key[19] , input \key[18] , input \key[17] , input \key[16] , input \key[15] , input \key[14] , input \key[13] , input \key[12] , input \key[11] , input \key[10] , input \key[9] , input \key[8] , input \key[7] , input \key[6] , input \key[5] , input \key[4] , input \key[3] , input \key[2] , input \key[1] , input \key[0] , input clk, output \data[19] , output \data[20] , output \data[21] , output \data[23] , output \data[24] , output \data[25] , output \data[26] , output \data[27] , output \data[28] , output \data[29] , output \data[30] , output \data[31] );

reg \data[18] = 0 ;
assign \data[17]  = \data[18] ;
assign \data[14]  = \data[18] ;
assign \data[11]  = \data[18] ;
assign \data[10]  = \data[18] ;
assign \data[6]  = \data[18] ;
assign \data[2]  = \data[18] ;
assign \data[0]  = \data[18] ;
assign \data[22]  = \data[18] ;
// (0, 1, 'span4_vert_b_0')
// (0, 1, 'span4_vert_t_12')
// (0, 2, 'span4_vert_b_12')
// (0, 3, 'io_0/D_OUT_0')
// (0, 3, 'io_0/PAD')
// (0, 3, 'io_1/D_OUT_0')
// (0, 3, 'io_1/PAD')
// (0, 3, 'local_g0_0')
// (0, 3, 'local_g1_0')
// (0, 3, 'span4_vert_b_8')
// (0, 4, 'span4_vert_b_4')
// (0, 5, 'io_0/D_OUT_0')
// (0, 5, 'io_0/PAD')
// (0, 5, 'local_g0_0')
// (0, 5, 'span4_horz_0')
// (0, 5, 'span4_horz_1')
// (0, 5, 'span4_vert_b_0')
// (0, 5, 'span4_vert_t_12')
// (0, 6, 'io_1/D_OUT_0')
// (0, 6, 'io_1/PAD')
// (0, 6, 'local_g1_4')
// (0, 6, 'span4_vert_b_12')
// (0, 7, 'io_0/D_OUT_0')
// (0, 7, 'io_0/PAD')
// (0, 7, 'local_g0_0')
// (0, 7, 'span4_vert_b_8')
// (0, 8, 'span4_vert_b_4')
// (0, 9, 'io_0/D_OUT_0')
// (0, 9, 'io_0/PAD')
// (0, 9, 'local_g1_1')
// (0, 9, 'span12_horz_1')
// (0, 9, 'span4_horz_0')
// (0, 9, 'span4_vert_b_0')
// (0, 9, 'span4_vert_t_12')
// (0, 10, 'span4_vert_b_12')
// (0, 11, 'io_0/D_OUT_0')
// (0, 11, 'io_0/PAD')
// (0, 11, 'local_g0_0')
// (0, 11, 'span4_vert_b_8')
// (0, 12, 'io_0/D_OUT_0')
// (0, 12, 'io_0/PAD')
// (0, 12, 'local_g0_4')
// (0, 12, 'span4_vert_b_4')
// (0, 13, 'span4_vert_b_0')
// (0, 20, 'logic_op_tnr_5')
// (0, 21, 'logic_op_rgt_5')
// (0, 21, 'span12_horz_1')
// (0, 22, 'logic_op_bnr_5')
// (1, 0, 'span4_horz_r_4')
// (1, 5, 'sp4_h_r_12')
// (1, 5, 'sp4_h_r_13')
// (1, 9, 'sp12_h_r_2')
// (1, 9, 'sp4_h_r_13')
// (1, 20, 'neigh_op_top_5')
// (1, 21, 'lutff_5/out')
// (1, 21, 'sp12_h_r_2')
// (1, 22, 'neigh_op_bot_5')
// (2, 0, 'span4_horz_r_8')
// (2, 5, 'sp4_h_r_24')
// (2, 5, 'sp4_h_r_25')
// (2, 9, 'sp12_h_r_5')
// (2, 9, 'sp4_h_r_24')
// (2, 20, 'neigh_op_tnl_5')
// (2, 21, 'neigh_op_lft_5')
// (2, 21, 'sp12_h_r_5')
// (2, 22, 'neigh_op_bnl_5')
// (3, 0, 'io_1/D_OUT_0')
// (3, 0, 'io_1/PAD')
// (3, 0, 'local_g1_4')
// (3, 0, 'span4_horz_r_12')
// (3, 2, 'sp4_r_v_b_45')
// (3, 3, 'sp4_r_v_b_32')
// (3, 4, 'sp4_r_v_b_21')
// (3, 5, 'sp4_h_r_36')
// (3, 5, 'sp4_h_r_37')
// (3, 5, 'sp4_r_v_b_8')
// (3, 6, 'sp4_r_v_b_37')
// (3, 7, 'sp4_r_v_b_24')
// (3, 8, 'sp4_r_v_b_13')
// (3, 9, 'sp12_h_r_6')
// (3, 9, 'sp4_h_r_37')
// (3, 9, 'sp4_r_v_b_0')
// (3, 21, 'sp12_h_r_6')
// (4, 0, 'span4_horz_l_12')
// (4, 1, 'sp4_v_t_45')
// (4, 2, 'sp4_v_b_45')
// (4, 3, 'sp4_v_b_32')
// (4, 4, 'sp4_v_b_21')
// (4, 5, 'sp4_h_l_36')
// (4, 5, 'sp4_h_l_37')
// (4, 5, 'sp4_v_b_8')
// (4, 5, 'sp4_v_t_37')
// (4, 6, 'sp4_v_b_37')
// (4, 7, 'sp4_v_b_24')
// (4, 8, 'sp4_v_b_13')
// (4, 9, 'sp12_h_r_9')
// (4, 9, 'sp4_h_l_37')
// (4, 9, 'sp4_v_b_0')
// (4, 21, 'sp12_h_r_9')
// (5, 9, 'sp12_h_r_10')
// (5, 21, 'sp12_h_r_10')
// (6, 9, 'sp12_h_r_13')
// (6, 21, 'sp12_h_r_13')
// (7, 9, 'sp12_h_r_14')
// (7, 21, 'sp12_h_r_14')
// (8, 9, 'sp12_h_r_17')
// (8, 21, 'sp12_h_r_17')
// (9, 9, 'sp12_h_r_18')
// (9, 21, 'sp12_h_r_18')
// (10, 9, 'sp12_h_r_21')
// (10, 21, 'sp12_h_r_21')
// (11, 9, 'sp12_h_r_22')
// (11, 21, 'sp12_h_r_22')
// (12, 9, 'sp12_h_l_22')
// (12, 9, 'sp12_v_t_22')
// (12, 10, 'sp12_v_b_22')
// (12, 11, 'sp12_v_b_21')
// (12, 12, 'sp12_v_b_18')
// (12, 13, 'sp12_v_b_17')
// (12, 14, 'sp12_v_b_14')
// (12, 15, 'sp12_v_b_13')
// (12, 16, 'sp12_v_b_10')
// (12, 17, 'sp12_v_b_9')
// (12, 18, 'sp12_v_b_6')
// (12, 19, 'sp12_v_b_5')
// (12, 20, 'sp12_v_b_2')
// (12, 21, 'sp12_h_l_22')
// (12, 21, 'sp12_v_b_1')

wire \data[16] ;
// (0, 4, 'io_0/D_OUT_0')
// (0, 4, 'io_0/PAD')

wire \data[15] ;
// (0, 4, 'io_1/D_OUT_0')
// (0, 4, 'io_1/PAD')

wire \data[13] ;
// (0, 5, 'io_1/D_OUT_0')
// (0, 5, 'io_1/PAD')

wire \data[12] ;
// (0, 6, 'io_0/D_OUT_0')
// (0, 6, 'io_0/PAD')

wire \data[9] ;
// (0, 7, 'io_1/D_OUT_0')
// (0, 7, 'io_1/PAD')

wire \data[8] ;
// (0, 8, 'io_0/D_OUT_0')
// (0, 8, 'io_0/PAD')

wire \data[7] ;
// (0, 8, 'io_1/D_OUT_0')
// (0, 8, 'io_1/PAD')

wire \data[5] ;
// (0, 9, 'io_1/D_OUT_0')
// (0, 9, 'io_1/PAD')

wire \data[4] ;
// (0, 10, 'io_0/D_OUT_0')
// (0, 10, 'io_0/PAD')

wire \data[3] ;
// (0, 10, 'io_1/D_OUT_0')
// (0, 10, 'io_1/PAD')

wire \data[1] ;
// (0, 11, 'io_1/D_OUT_0')
// (0, 11, 'io_1/PAD')

wire \key[31] ;
// (0, 12, 'io_1/D_IN_0')
// (0, 12, 'io_1/PAD')
// (0, 12, 'span4_horz_28')
// (1, 11, 'neigh_op_tnl_2')
// (1, 11, 'neigh_op_tnl_6')
// (1, 12, 'neigh_op_lft_2')
// (1, 12, 'neigh_op_lft_6')
// (1, 12, 'sp4_h_r_41')
// (1, 13, 'neigh_op_bnl_2')
// (1, 13, 'neigh_op_bnl_6')
// (1, 13, 'sp4_r_v_b_41')
// (1, 14, 'local_g1_4')
// (1, 14, 'lutff_6/in_3')
// (1, 14, 'sp4_r_v_b_28')
// (1, 15, 'sp4_r_v_b_17')
// (1, 16, 'sp4_r_v_b_4')
// (2, 12, 'sp4_h_l_41')
// (2, 12, 'sp4_v_t_41')
// (2, 13, 'sp4_v_b_41')
// (2, 14, 'sp4_v_b_28')
// (2, 15, 'sp4_v_b_17')
// (2, 16, 'sp4_v_b_4')

wire \key[30] ;
// (0, 12, 'span4_vert_t_12')
// (0, 13, 'io_0/D_IN_0')
// (0, 13, 'io_0/PAD')
// (0, 13, 'span4_vert_b_12')
// (0, 14, 'span4_vert_b_8')
// (0, 15, 'span4_vert_b_4')
// (0, 16, 'span4_horz_1')
// (0, 16, 'span4_vert_b_0')
// (1, 12, 'neigh_op_tnl_0')
// (1, 12, 'neigh_op_tnl_4')
// (1, 13, 'neigh_op_lft_0')
// (1, 13, 'neigh_op_lft_4')
// (1, 14, 'neigh_op_bnl_0')
// (1, 14, 'neigh_op_bnl_4')
// (1, 16, 'local_g0_4')
// (1, 16, 'lutff_1/in_3')
// (1, 16, 'sp4_h_r_12')
// (2, 16, 'sp4_h_r_25')
// (3, 16, 'sp4_h_r_36')
// (4, 16, 'sp4_h_l_36')

wire \key[29] ;
// (0, 13, 'io_1/D_IN_0')
// (0, 13, 'io_1/PAD')
// (0, 13, 'span4_horz_44')
// (1, 12, 'neigh_op_tnl_2')
// (1, 12, 'neigh_op_tnl_6')
// (1, 13, 'neigh_op_lft_2')
// (1, 13, 'neigh_op_lft_6')
// (1, 13, 'sp4_h_l_44')
// (1, 13, 'sp4_v_t_39')
// (1, 14, 'neigh_op_bnl_2')
// (1, 14, 'neigh_op_bnl_6')
// (1, 14, 'sp4_v_b_39')
// (1, 15, 'sp4_v_b_26')
// (1, 16, 'local_g0_7')
// (1, 16, 'lutff_1/in_2')
// (1, 16, 'sp4_v_b_15')
// (1, 17, 'sp4_v_b_2')

wire n16;
// (0, 13, 'logic_op_tnr_6')
// (0, 14, 'logic_op_rgt_6')
// (0, 15, 'logic_op_bnr_6')
// (1, 13, 'neigh_op_top_6')
// (1, 13, 'sp4_v_t_44')
// (1, 14, 'lutff_6/out')
// (1, 14, 'sp4_v_b_44')
// (1, 15, 'neigh_op_bot_6')
// (1, 15, 'sp4_v_b_33')
// (1, 16, 'sp4_v_b_20')
// (1, 17, 'sp4_v_b_9')
// (1, 17, 'sp4_v_t_37')
// (1, 18, 'sp4_v_b_37')
// (1, 19, 'sp4_v_b_24')
// (1, 20, 'sp4_v_b_13')
// (1, 21, 'local_g0_0')
// (1, 21, 'lutff_4/in_2')
// (1, 21, 'sp4_v_b_0')
// (2, 13, 'neigh_op_tnl_6')
// (2, 14, 'neigh_op_lft_6')
// (2, 15, 'neigh_op_bnl_6')

wire \key[28] ;
// (0, 14, 'io_0/D_IN_0')
// (0, 14, 'io_0/PAD')
// (1, 13, 'neigh_op_tnl_0')
// (1, 13, 'neigh_op_tnl_4')
// (1, 14, 'local_g0_4')
// (1, 14, 'lutff_6/in_2')
// (1, 14, 'neigh_op_lft_0')
// (1, 14, 'neigh_op_lft_4')
// (1, 15, 'neigh_op_bnl_0')
// (1, 15, 'neigh_op_bnl_4')

wire \key[27] ;
// (0, 14, 'io_1/D_IN_0')
// (0, 14, 'io_1/PAD')
// (1, 13, 'neigh_op_tnl_2')
// (1, 13, 'neigh_op_tnl_6')
// (1, 14, 'local_g1_2')
// (1, 14, 'lutff_6/in_1')
// (1, 14, 'neigh_op_lft_2')
// (1, 14, 'neigh_op_lft_6')
// (1, 15, 'neigh_op_bnl_2')
// (1, 15, 'neigh_op_bnl_6')

wire n19;
// (0, 15, 'logic_op_tnr_1')
// (0, 16, 'logic_op_rgt_1')
// (0, 17, 'logic_op_bnr_1')
// (1, 13, 'sp12_v_t_22')
// (1, 14, 'sp12_v_b_22')
// (1, 15, 'neigh_op_top_1')
// (1, 15, 'sp12_v_b_21')
// (1, 16, 'lutff_1/out')
// (1, 16, 'sp12_v_b_18')
// (1, 17, 'neigh_op_bot_1')
// (1, 17, 'sp12_v_b_17')
// (1, 18, 'sp12_v_b_14')
// (1, 19, 'sp12_v_b_13')
// (1, 20, 'sp12_v_b_10')
// (1, 21, 'sp12_v_b_9')
// (1, 22, 'local_g2_6')
// (1, 22, 'lutff_3/in_3')
// (1, 22, 'sp12_v_b_6')
// (1, 23, 'sp12_v_b_5')
// (1, 24, 'sp12_v_b_2')
// (1, 25, 'sp12_v_b_1')
// (2, 15, 'neigh_op_tnl_1')
// (2, 16, 'neigh_op_lft_1')
// (2, 17, 'neigh_op_bnl_1')

wire \key[26] ;
// (0, 16, 'io_0/D_IN_0')
// (0, 16, 'io_0/PAD')
// (0, 16, 'span4_horz_24')
// (1, 13, 'sp4_r_v_b_37')
// (1, 14, 'local_g0_0')
// (1, 14, 'lutff_6/in_0')
// (1, 14, 'sp4_r_v_b_24')
// (1, 15, 'neigh_op_tnl_0')
// (1, 15, 'neigh_op_tnl_4')
// (1, 15, 'sp4_r_v_b_13')
// (1, 16, 'neigh_op_lft_0')
// (1, 16, 'neigh_op_lft_4')
// (1, 16, 'sp4_h_r_37')
// (1, 16, 'sp4_r_v_b_0')
// (1, 17, 'neigh_op_bnl_0')
// (1, 17, 'neigh_op_bnl_4')
// (2, 12, 'sp4_v_t_37')
// (2, 13, 'sp4_v_b_37')
// (2, 14, 'sp4_v_b_24')
// (2, 15, 'sp4_v_b_13')
// (2, 16, 'sp4_h_l_37')
// (2, 16, 'sp4_v_b_0')

wire \key[25] ;
// (0, 16, 'io_1/D_IN_0')
// (0, 16, 'io_1/PAD')
// (1, 15, 'neigh_op_tnl_2')
// (1, 15, 'neigh_op_tnl_6')
// (1, 16, 'local_g0_2')
// (1, 16, 'lutff_1/in_1')
// (1, 16, 'neigh_op_lft_2')
// (1, 16, 'neigh_op_lft_6')
// (1, 17, 'neigh_op_bnl_2')
// (1, 17, 'neigh_op_bnl_6')

wire \key[24] ;
// (0, 17, 'io_0/D_IN_0')
// (0, 17, 'io_0/PAD')
// (1, 16, 'neigh_op_tnl_0')
// (1, 16, 'neigh_op_tnl_4')
// (1, 17, 'neigh_op_lft_0')
// (1, 17, 'neigh_op_lft_4')
// (1, 18, 'local_g2_0')
// (1, 18, 'lutff_5/in_3')
// (1, 18, 'neigh_op_bnl_0')
// (1, 18, 'neigh_op_bnl_4')

wire \key[23] ;
// (0, 17, 'io_1/D_IN_0')
// (0, 17, 'io_1/PAD')
// (1, 16, 'neigh_op_tnl_2')
// (1, 16, 'neigh_op_tnl_6')
// (1, 17, 'neigh_op_lft_2')
// (1, 17, 'neigh_op_lft_6')
// (1, 18, 'local_g3_2')
// (1, 18, 'lutff_5/in_2')
// (1, 18, 'neigh_op_bnl_2')
// (1, 18, 'neigh_op_bnl_6')

wire n24;
// (0, 17, 'logic_op_tnr_5')
// (0, 18, 'logic_op_rgt_5')
// (0, 19, 'logic_op_bnr_5')
// (1, 17, 'neigh_op_top_5')
// (1, 17, 'sp4_v_t_42')
// (1, 18, 'lutff_5/out')
// (1, 18, 'sp4_v_b_42')
// (1, 19, 'neigh_op_bot_5')
// (1, 19, 'sp4_v_b_31')
// (1, 20, 'sp4_v_b_18')
// (1, 21, 'local_g0_7')
// (1, 21, 'lutff_4/in_3')
// (1, 21, 'sp4_v_b_7')
// (2, 17, 'neigh_op_tnl_5')
// (2, 18, 'neigh_op_lft_5')
// (2, 19, 'neigh_op_bnl_5')

wire \key[22] ;
// (0, 18, 'io_0/D_IN_0')
// (0, 18, 'io_0/PAD')
// (0, 18, 'span4_horz_32')
// (1, 15, 'sp4_r_v_b_45')
// (1, 16, 'local_g0_3')
// (1, 16, 'lutff_1/in_0')
// (1, 16, 'sp4_r_v_b_32')
// (1, 17, 'neigh_op_tnl_0')
// (1, 17, 'neigh_op_tnl_4')
// (1, 17, 'sp4_r_v_b_21')
// (1, 18, 'neigh_op_lft_0')
// (1, 18, 'neigh_op_lft_4')
// (1, 18, 'sp4_h_r_45')
// (1, 18, 'sp4_r_v_b_8')
// (1, 19, 'neigh_op_bnl_0')
// (1, 19, 'neigh_op_bnl_4')
// (2, 14, 'sp4_v_t_45')
// (2, 15, 'sp4_v_b_45')
// (2, 16, 'sp4_v_b_32')
// (2, 17, 'sp4_v_b_21')
// (2, 18, 'sp4_h_l_45')
// (2, 18, 'sp4_v_b_8')

wire \key[21] ;
// (0, 18, 'io_1/D_IN_0')
// (0, 18, 'io_1/PAD')
// (1, 17, 'neigh_op_tnl_2')
// (1, 17, 'neigh_op_tnl_6')
// (1, 18, 'local_g0_2')
// (1, 18, 'lutff_5/in_1')
// (1, 18, 'neigh_op_lft_2')
// (1, 18, 'neigh_op_lft_6')
// (1, 19, 'neigh_op_bnl_2')
// (1, 19, 'neigh_op_bnl_6')

wire \key[20] ;
// (0, 18, 'span4_vert_t_12')
// (0, 19, 'io_0/D_IN_0')
// (0, 19, 'io_0/PAD')
// (0, 19, 'span4_vert_b_12')
// (0, 20, 'span4_vert_b_8')
// (0, 21, 'span4_vert_b_4')
// (0, 22, 'span4_horz_1')
// (0, 22, 'span4_vert_b_0')
// (1, 18, 'neigh_op_tnl_0')
// (1, 18, 'neigh_op_tnl_4')
// (1, 19, 'neigh_op_lft_0')
// (1, 19, 'neigh_op_lft_4')
// (1, 20, 'neigh_op_bnl_0')
// (1, 20, 'neigh_op_bnl_4')
// (1, 22, 'local_g0_4')
// (1, 22, 'lutff_7/in_3')
// (1, 22, 'sp4_h_r_12')
// (2, 22, 'sp4_h_r_25')
// (3, 22, 'sp4_h_r_36')
// (4, 22, 'sp4_h_l_36')

wire \key[19] ;
// (0, 19, 'io_1/D_IN_0')
// (0, 19, 'io_1/PAD')
// (0, 19, 'span4_horz_36')
// (1, 18, 'neigh_op_tnl_2')
// (1, 18, 'neigh_op_tnl_6')
// (1, 19, 'neigh_op_lft_2')
// (1, 19, 'neigh_op_lft_6')
// (1, 19, 'sp4_h_l_36')
// (1, 19, 'sp4_v_t_43')
// (1, 20, 'neigh_op_bnl_2')
// (1, 20, 'neigh_op_bnl_6')
// (1, 20, 'sp4_v_b_43')
// (1, 21, 'sp4_v_b_30')
// (1, 22, 'local_g0_3')
// (1, 22, 'lutff_7/in_2')
// (1, 22, 'sp4_v_b_19')
// (1, 23, 'sp4_v_b_6')

wire \key[18] ;
// (0, 20, 'io_0/D_IN_0')
// (0, 20, 'io_0/PAD')
// (0, 20, 'span4_horz_32')
// (1, 17, 'sp4_r_v_b_45')
// (1, 18, 'local_g0_3')
// (1, 18, 'lutff_5/in_0')
// (1, 18, 'sp4_r_v_b_32')
// (1, 19, 'neigh_op_tnl_0')
// (1, 19, 'neigh_op_tnl_4')
// (1, 19, 'sp4_r_v_b_21')
// (1, 20, 'neigh_op_lft_0')
// (1, 20, 'neigh_op_lft_4')
// (1, 20, 'sp4_h_r_45')
// (1, 20, 'sp4_r_v_b_8')
// (1, 21, 'neigh_op_bnl_0')
// (1, 21, 'neigh_op_bnl_4')
// (2, 16, 'sp4_v_t_45')
// (2, 17, 'sp4_v_b_45')
// (2, 18, 'sp4_v_b_32')
// (2, 19, 'sp4_v_b_21')
// (2, 20, 'sp4_h_l_45')
// (2, 20, 'sp4_v_b_8')

wire \key[17] ;
// (0, 20, 'io_1/D_IN_0')
// (0, 20, 'io_1/PAD')
// (1, 19, 'neigh_op_tnl_2')
// (1, 19, 'neigh_op_tnl_6')
// (1, 20, 'neigh_op_lft_2')
// (1, 20, 'neigh_op_lft_6')
// (1, 21, 'local_g2_6')
// (1, 21, 'lutff_3/in_3')
// (1, 21, 'neigh_op_bnl_2')
// (1, 21, 'neigh_op_bnl_6')

wire n31;
// (0, 20, 'logic_op_tnr_3')
// (0, 21, 'logic_op_rgt_3')
// (0, 22, 'logic_op_bnr_3')
// (1, 20, 'neigh_op_top_3')
// (1, 21, 'local_g1_3')
// (1, 21, 'lutff_3/out')
// (1, 21, 'lutff_4/in_0')
// (1, 22, 'neigh_op_bot_3')
// (2, 20, 'neigh_op_tnl_3')
// (2, 21, 'neigh_op_lft_3')
// (2, 22, 'neigh_op_bnl_3')

wire n32;
// (0, 20, 'logic_op_tnr_4')
// (0, 21, 'logic_op_rgt_4')
// (0, 22, 'logic_op_bnr_4')
// (1, 20, 'neigh_op_top_4')
// (1, 21, 'local_g1_4')
// (1, 21, 'lutff_4/out')
// (1, 21, 'lutff_5/in_0')
// (1, 22, 'neigh_op_bot_4')
// (2, 20, 'neigh_op_tnl_4')
// (2, 21, 'neigh_op_lft_4')
// (2, 22, 'neigh_op_bnl_4')

wire \key[16] ;
// (0, 21, 'io_0/D_IN_0')
// (0, 21, 'io_0/PAD')
// (0, 21, 'span12_horz_0')
// (1, 20, 'neigh_op_tnl_0')
// (1, 20, 'neigh_op_tnl_4')
// (1, 21, 'local_g0_3')
// (1, 21, 'lutff_3/in_2')
// (1, 21, 'neigh_op_lft_0')
// (1, 21, 'neigh_op_lft_4')
// (1, 21, 'sp12_h_r_3')
// (1, 22, 'neigh_op_bnl_0')
// (1, 22, 'neigh_op_bnl_4')
// (2, 21, 'sp12_h_r_4')
// (3, 21, 'sp12_h_r_7')
// (4, 21, 'sp12_h_r_8')
// (5, 21, 'sp12_h_r_11')
// (6, 21, 'sp12_h_r_12')
// (7, 21, 'sp12_h_r_15')
// (8, 21, 'sp12_h_r_16')
// (9, 21, 'sp12_h_r_19')
// (10, 21, 'sp12_h_r_20')
// (11, 21, 'sp12_h_r_23')
// (12, 21, 'sp12_h_l_23')

wire \key[15] ;
// (0, 21, 'io_1/D_IN_0')
// (0, 21, 'io_1/PAD')
// (1, 20, 'neigh_op_tnl_2')
// (1, 20, 'neigh_op_tnl_6')
// (1, 21, 'local_g0_2')
// (1, 21, 'lutff_3/in_1')
// (1, 21, 'neigh_op_lft_2')
// (1, 21, 'neigh_op_lft_6')
// (1, 22, 'neigh_op_bnl_2')
// (1, 22, 'neigh_op_bnl_6')

wire n35;
// (0, 21, 'logic_op_tnr_3')
// (0, 22, 'logic_op_rgt_3')
// (0, 23, 'logic_op_bnr_3')
// (1, 20, 'sp4_r_v_b_47')
// (1, 21, 'local_g2_2')
// (1, 21, 'lutff_5/in_1')
// (1, 21, 'neigh_op_top_3')
// (1, 21, 'sp4_r_v_b_34')
// (1, 22, 'lutff_3/out')
// (1, 22, 'sp4_r_v_b_23')
// (1, 23, 'neigh_op_bot_3')
// (1, 23, 'sp4_r_v_b_10')
// (2, 19, 'sp4_v_t_47')
// (2, 20, 'sp4_v_b_47')
// (2, 21, 'neigh_op_tnl_3')
// (2, 21, 'sp4_v_b_34')
// (2, 22, 'neigh_op_lft_3')
// (2, 22, 'sp4_v_b_23')
// (2, 23, 'neigh_op_bnl_3')
// (2, 23, 'sp4_v_b_10')

wire n36;
// (0, 21, 'logic_op_tnr_7')
// (0, 22, 'logic_op_rgt_7')
// (0, 23, 'logic_op_bnr_7')
// (1, 21, 'neigh_op_top_7')
// (1, 22, 'local_g0_7')
// (1, 22, 'lutff_3/in_0')
// (1, 22, 'lutff_7/out')
// (1, 23, 'neigh_op_bot_7')
// (2, 21, 'neigh_op_tnl_7')
// (2, 22, 'neigh_op_lft_7')
// (2, 23, 'neigh_op_bnl_7')

wire \key[14] ;
// (0, 22, 'io_0/D_IN_0')
// (0, 22, 'io_0/PAD')
// (1, 21, 'neigh_op_tnl_0')
// (1, 21, 'neigh_op_tnl_4')
// (1, 22, 'local_g0_0')
// (1, 22, 'lutff_7/in_1')
// (1, 22, 'neigh_op_lft_0')
// (1, 22, 'neigh_op_lft_4')
// (1, 23, 'neigh_op_bnl_0')
// (1, 23, 'neigh_op_bnl_4')

wire \key[13] ;
// (0, 22, 'io_1/D_IN_0')
// (0, 22, 'io_1/PAD')
// (1, 21, 'neigh_op_tnl_2')
// (1, 21, 'neigh_op_tnl_6')
// (1, 22, 'local_g1_2')
// (1, 22, 'lutff_7/in_0')
// (1, 22, 'neigh_op_lft_2')
// (1, 22, 'neigh_op_lft_6')
// (1, 23, 'neigh_op_bnl_2')
// (1, 23, 'neigh_op_bnl_6')

wire \key[12] ;
// (0, 23, 'io_0/D_IN_0')
// (0, 23, 'io_0/PAD')
// (0, 23, 'span4_horz_24')
// (1, 20, 'sp4_r_v_b_37')
// (1, 21, 'local_g1_0')
// (1, 21, 'lutff_3/in_0')
// (1, 21, 'sp4_r_v_b_24')
// (1, 22, 'neigh_op_tnl_0')
// (1, 22, 'neigh_op_tnl_4')
// (1, 22, 'sp4_r_v_b_13')
// (1, 23, 'neigh_op_lft_0')
// (1, 23, 'neigh_op_lft_4')
// (1, 23, 'sp4_h_r_37')
// (1, 23, 'sp4_r_v_b_0')
// (1, 24, 'neigh_op_bnl_0')
// (1, 24, 'neigh_op_bnl_4')
// (2, 19, 'sp4_v_t_37')
// (2, 20, 'sp4_v_b_37')
// (2, 21, 'sp4_v_b_24')
// (2, 22, 'sp4_v_b_13')
// (2, 23, 'sp4_h_l_37')
// (2, 23, 'sp4_v_b_0')

wire \key[11] ;
// (0, 23, 'io_1/D_IN_0')
// (0, 23, 'io_1/PAD')
// (1, 22, 'neigh_op_tnl_2')
// (1, 22, 'neigh_op_tnl_6')
// (1, 23, 'neigh_op_lft_2')
// (1, 23, 'neigh_op_lft_6')
// (1, 24, 'local_g3_2')
// (1, 24, 'lutff_2/in_3')
// (1, 24, 'neigh_op_bnl_2')
// (1, 24, 'neigh_op_bnl_6')

wire n41;
// (0, 23, 'logic_op_tnr_2')
// (0, 24, 'logic_op_rgt_2')
// (0, 25, 'logic_op_bnr_2')
// (1, 20, 'sp4_v_t_41')
// (1, 21, 'local_g2_1')
// (1, 21, 'lutff_4/in_1')
// (1, 21, 'sp4_v_b_41')
// (1, 22, 'sp4_v_b_28')
// (1, 23, 'neigh_op_top_2')
// (1, 23, 'sp4_v_b_17')
// (1, 24, 'lutff_2/out')
// (1, 24, 'sp4_v_b_4')
// (1, 25, 'neigh_op_bot_2')
// (2, 23, 'neigh_op_tnl_2')
// (2, 24, 'neigh_op_lft_2')
// (2, 25, 'neigh_op_bnl_2')

wire \key[10] ;
// (0, 24, 'io_0/D_IN_0')
// (0, 24, 'io_0/PAD')
// (1, 23, 'neigh_op_tnl_0')
// (1, 23, 'neigh_op_tnl_4')
// (1, 24, 'local_g0_0')
// (1, 24, 'lutff_2/in_2')
// (1, 24, 'neigh_op_lft_0')
// (1, 24, 'neigh_op_lft_4')
// (1, 25, 'neigh_op_bnl_0')
// (1, 25, 'neigh_op_bnl_4')

wire \key[9] ;
// (0, 24, 'io_1/D_IN_0')
// (0, 24, 'io_1/PAD')
// (1, 23, 'neigh_op_tnl_2')
// (1, 23, 'neigh_op_tnl_6')
// (1, 24, 'local_g1_2')
// (1, 24, 'lutff_2/in_1')
// (1, 24, 'neigh_op_lft_2')
// (1, 24, 'neigh_op_lft_6')
// (1, 25, 'neigh_op_bnl_2')
// (1, 25, 'neigh_op_bnl_6')

wire \key[8] ;
// (0, 25, 'io_0/D_IN_0')
// (0, 25, 'io_0/PAD')
// (1, 24, 'local_g2_0')
// (1, 24, 'lutff_2/in_0')
// (1, 24, 'neigh_op_tnl_0')
// (1, 24, 'neigh_op_tnl_4')
// (1, 25, 'neigh_op_lft_0')
// (1, 25, 'neigh_op_lft_4')
// (1, 26, 'neigh_op_bnl_0')
// (1, 26, 'neigh_op_bnl_4')

wire \key[7] ;
// (0, 25, 'io_1/D_IN_0')
// (0, 25, 'io_1/PAD')
// (0, 25, 'span4_horz_28')
// (1, 24, 'neigh_op_tnl_2')
// (1, 24, 'neigh_op_tnl_6')
// (1, 25, 'neigh_op_lft_2')
// (1, 25, 'neigh_op_lft_6')
// (1, 25, 'sp4_h_r_41')
// (1, 26, 'neigh_op_bnl_2')
// (1, 26, 'neigh_op_bnl_6')
// (1, 26, 'sp4_r_v_b_41')
// (1, 27, 'local_g1_4')
// (1, 27, 'lutff_4/in_3')
// (1, 27, 'sp4_r_v_b_28')
// (1, 28, 'sp4_r_v_b_17')
// (1, 29, 'sp4_r_v_b_4')
// (2, 25, 'sp4_h_l_41')
// (2, 25, 'sp4_v_t_41')
// (2, 26, 'sp4_v_b_41')
// (2, 27, 'sp4_v_b_28')
// (2, 28, 'sp4_v_b_17')
// (2, 29, 'sp4_v_b_4')

wire n46;
// (0, 26, 'logic_op_tnr_4')
// (0, 27, 'logic_op_rgt_4')
// (0, 28, 'logic_op_bnr_4')
// (1, 19, 'sp12_v_t_23')
// (1, 20, 'sp12_v_b_23')
// (1, 21, 'sp12_v_b_20')
// (1, 22, 'local_g2_3')
// (1, 22, 'lutff_3/in_2')
// (1, 22, 'sp12_v_b_19')
// (1, 23, 'sp12_v_b_16')
// (1, 24, 'sp12_v_b_15')
// (1, 25, 'sp12_v_b_12')
// (1, 26, 'neigh_op_top_4')
// (1, 26, 'sp12_v_b_11')
// (1, 27, 'lutff_4/out')
// (1, 27, 'sp12_v_b_8')
// (1, 28, 'neigh_op_bot_4')
// (1, 28, 'sp12_v_b_7')
// (1, 29, 'sp12_v_b_4')
// (1, 30, 'sp12_v_b_3')
// (1, 31, 'sp12_v_b_0')
// (2, 26, 'neigh_op_tnl_4')
// (2, 27, 'neigh_op_lft_4')
// (2, 28, 'neigh_op_bnl_4')

wire \key[6] ;
// (0, 27, 'io_0/D_IN_0')
// (0, 27, 'io_0/PAD')
// (1, 26, 'neigh_op_tnl_0')
// (1, 26, 'neigh_op_tnl_4')
// (1, 27, 'local_g0_0')
// (1, 27, 'lutff_4/in_2')
// (1, 27, 'neigh_op_lft_0')
// (1, 27, 'neigh_op_lft_4')
// (1, 28, 'neigh_op_bnl_0')
// (1, 28, 'neigh_op_bnl_4')

wire \key[5] ;
// (0, 27, 'io_1/D_IN_0')
// (0, 27, 'io_1/PAD')
// (1, 26, 'neigh_op_tnl_2')
// (1, 26, 'neigh_op_tnl_6')
// (1, 27, 'local_g1_2')
// (1, 27, 'lutff_4/in_1')
// (1, 27, 'neigh_op_lft_2')
// (1, 27, 'neigh_op_lft_6')
// (1, 28, 'neigh_op_bnl_2')
// (1, 28, 'neigh_op_bnl_6')

wire \key[4] ;
// (0, 28, 'io_0/D_IN_0')
// (0, 28, 'io_0/PAD')
// (1, 27, 'local_g2_0')
// (1, 27, 'lutff_4/in_0')
// (1, 27, 'neigh_op_tnl_0')
// (1, 27, 'neigh_op_tnl_4')
// (1, 28, 'neigh_op_lft_0')
// (1, 28, 'neigh_op_lft_4')
// (1, 29, 'neigh_op_bnl_0')
// (1, 29, 'neigh_op_bnl_4')

wire \key[3] ;
// (0, 28, 'io_1/D_IN_0')
// (0, 28, 'io_1/PAD')
// (0, 28, 'span4_horz_28')
// (1, 27, 'neigh_op_tnl_2')
// (1, 27, 'neigh_op_tnl_6')
// (1, 28, 'neigh_op_lft_2')
// (1, 28, 'neigh_op_lft_6')
// (1, 28, 'sp4_h_r_41')
// (1, 29, 'neigh_op_bnl_2')
// (1, 29, 'neigh_op_bnl_6')
// (1, 29, 'sp4_r_v_b_41')
// (1, 30, 'local_g0_4')
// (1, 30, 'lutff_1/in_3')
// (1, 30, 'sp4_r_v_b_28')
// (1, 31, 'sp4_r_v_b_17')
// (1, 32, 'sp4_r_v_b_4')
// (2, 28, 'sp4_h_l_41')
// (2, 28, 'sp4_v_t_41')
// (2, 29, 'sp4_v_b_41')
// (2, 30, 'sp4_v_b_28')
// (2, 31, 'sp4_v_b_17')
// (2, 32, 'sp4_v_b_4')

wire n51;
// (0, 29, 'logic_op_tnr_1')
// (0, 30, 'logic_op_rgt_1')
// (0, 31, 'logic_op_bnr_1')
// (1, 19, 'sp12_v_t_22')
// (1, 20, 'sp12_v_b_22')
// (1, 21, 'sp12_v_b_21')
// (1, 22, 'local_g2_2')
// (1, 22, 'lutff_3/in_1')
// (1, 22, 'sp12_v_b_18')
// (1, 23, 'sp12_v_b_17')
// (1, 24, 'sp12_v_b_14')
// (1, 25, 'sp12_v_b_13')
// (1, 26, 'sp12_v_b_10')
// (1, 27, 'sp12_v_b_9')
// (1, 28, 'sp12_v_b_6')
// (1, 29, 'neigh_op_top_1')
// (1, 29, 'sp12_v_b_5')
// (1, 30, 'lutff_1/out')
// (1, 30, 'sp12_v_b_2')
// (1, 31, 'neigh_op_bot_1')
// (1, 31, 'sp12_v_b_1')
// (2, 29, 'neigh_op_tnl_1')
// (2, 30, 'neigh_op_lft_1')
// (2, 31, 'neigh_op_bnl_1')

wire \key[2] ;
// (0, 30, 'io_0/D_IN_0')
// (0, 30, 'io_0/PAD')
// (1, 29, 'neigh_op_tnl_0')
// (1, 29, 'neigh_op_tnl_4')
// (1, 30, 'local_g1_0')
// (1, 30, 'lutff_1/in_2')
// (1, 30, 'neigh_op_lft_0')
// (1, 30, 'neigh_op_lft_4')
// (1, 31, 'neigh_op_bnl_0')
// (1, 31, 'neigh_op_bnl_4')

wire \key[1] ;
// (0, 30, 'io_1/D_IN_0')
// (0, 30, 'io_1/PAD')
// (1, 29, 'neigh_op_tnl_2')
// (1, 29, 'neigh_op_tnl_6')
// (1, 30, 'local_g0_2')
// (1, 30, 'lutff_1/in_1')
// (1, 30, 'neigh_op_lft_2')
// (1, 30, 'neigh_op_lft_6')
// (1, 31, 'neigh_op_bnl_2')
// (1, 31, 'neigh_op_bnl_6')

wire \key[0] ;
// (0, 31, 'io_0/D_IN_0')
// (0, 31, 'io_0/PAD')
// (1, 30, 'local_g3_0')
// (1, 30, 'lutff_1/in_0')
// (1, 30, 'neigh_op_tnl_0')
// (1, 30, 'neigh_op_tnl_4')
// (1, 31, 'neigh_op_lft_0')
// (1, 31, 'neigh_op_lft_4')
// (1, 32, 'neigh_op_bnl_0')
// (1, 32, 'neigh_op_bnl_4')

wire clk;
// (0, 31, 'io_1/D_IN_0')
// (0, 31, 'io_1/PAD')
// (0, 31, 'span12_horz_20')
// (1, 20, 'sp4_r_v_b_45')
// (1, 21, 'local_g2_0')
// (1, 21, 'lutff_global/clk')
// (1, 21, 'sp4_r_v_b_32')
// (1, 22, 'sp4_r_v_b_21')
// (1, 23, 'sp4_r_v_b_8')
// (1, 30, 'neigh_op_tnl_2')
// (1, 30, 'neigh_op_tnl_6')
// (1, 31, 'neigh_op_lft_2')
// (1, 31, 'neigh_op_lft_6')
// (1, 31, 'sp12_h_r_23')
// (1, 32, 'neigh_op_bnl_2')
// (1, 32, 'neigh_op_bnl_6')
// (2, 19, 'sp12_v_t_23')
// (2, 19, 'sp4_v_t_45')
// (2, 20, 'sp12_v_b_23')
// (2, 20, 'sp4_v_b_45')
// (2, 21, 'sp12_v_b_20')
// (2, 21, 'sp4_v_b_32')
// (2, 22, 'sp12_v_b_19')
// (2, 22, 'sp4_v_b_21')
// (2, 23, 'sp12_v_b_16')
// (2, 23, 'sp4_v_b_8')
// (2, 24, 'sp12_v_b_15')
// (2, 25, 'sp12_v_b_12')
// (2, 26, 'sp12_v_b_11')
// (2, 27, 'sp12_v_b_8')
// (2, 28, 'sp12_v_b_7')
// (2, 29, 'sp12_v_b_4')
// (2, 30, 'sp12_v_b_3')
// (2, 31, 'sp12_h_l_23')
// (2, 31, 'sp12_v_b_0')

wire \data[19] ;
// (2, 0, 'io_0/D_OUT_0')
// (2, 0, 'io_0/PAD')

wire \data[20] ;
// (2, 0, 'io_1/D_OUT_0')
// (2, 0, 'io_1/PAD')

wire \data[21] ;
// (3, 0, 'io_0/D_OUT_0')
// (3, 0, 'io_0/PAD')

wire \data[23] ;
// (4, 0, 'io_0/D_OUT_0')
// (4, 0, 'io_0/PAD')

wire \data[24] ;
// (4, 0, 'io_1/D_OUT_0')
// (4, 0, 'io_1/PAD')

wire \data[25] ;
// (5, 0, 'io_0/D_OUT_0')
// (5, 0, 'io_0/PAD')

wire \data[26] ;
// (5, 0, 'io_1/D_OUT_0')
// (5, 0, 'io_1/PAD')

wire \data[27] ;
// (6, 0, 'io_0/D_OUT_0')
// (6, 0, 'io_0/PAD')

wire \data[28] ;
// (6, 0, 'io_1/D_OUT_0')
// (6, 0, 'io_1/PAD')

wire \data[29] ;
// (7, 0, 'io_1/D_OUT_0')
// (7, 0, 'io_1/PAD')

wire \data[30] ;
// (8, 0, 'io_0/D_OUT_0')
// (8, 0, 'io_0/PAD')

wire \data[31] ;
// (9, 0, 'io_0/D_OUT_0')
// (9, 0, 'io_0/PAD')

wire n68;
// (1, 21, 'lutff_5/lout')

wire n69;
// (1, 18, 'lutff_5/lout')

wire n70;
// (1, 27, 'lutff_4/lout')

wire n71;
// (1, 14, 'lutff_6/lout')

wire n72;
// (1, 21, 'lutff_4/lout')

wire n73;
// (1, 24, 'lutff_2/lout')

wire n74;
// (1, 21, 'lutff_3/lout')

wire n75;
// (1, 30, 'lutff_1/lout')

wire n76;
// (1, 22, 'lutff_3/lout')

wire n77;
// (1, 22, 'lutff_7/lout')

wire n78;
// (1, 16, 'lutff_1/lout')

assign n68 = /* LUT    1 21  5 */ 1'b0 ? 1'b0 : 1'b0 ? 1'b0 : n35 ? n32 ? 1'b1 : 1'b0 : 1'b0;
assign n69 = /* LUT    1 18  5 */ \key[24]  ? \key[23]  ? \key[21]  ? \key[18]  ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n70 = /* LUT    1 27  4 */ \key[7]  ? \key[6]  ? \key[5]  ? \key[4]  ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n71 = /* LUT    1 14  6 */ \key[31]  ? \key[28]  ? \key[27]  ? \key[26]  ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n72 = /* LUT    1 21  4 */ n24 ? n16 ? n41 ? n31 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n73 = /* LUT    1 24  2 */ \key[11]  ? \key[10]  ? \key[9]  ? \key[8]  ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n74 = /* LUT    1 21  3 */ \key[17]  ? \key[16]  ? \key[15]  ? \key[12]  ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n75 = /* LUT    1 30  1 */ \key[3]  ? 1'b0 : \key[2]  ? 1'b0 : \key[1]  ? 1'b0 : \key[0]  ? 1'b0 : 1'b1;
assign n76 = /* LUT    1 22  3 */ n19 ? n46 ? n51 ? n36 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n77 = /* LUT    1 22  7 */ \key[20]  ? 1'b0 : \key[19]  ? 1'b0 : \key[14]  ? 1'b0 : \key[13]  ? 1'b0 : 1'b1;
assign n78 = /* LUT    1 16  1 */ \key[30]  ? 1'b0 : \key[29]  ? 1'b0 : \key[25]  ? 1'b0 : \key[22]  ? 1'b0 : 1'b1;
/* FF  1 21  5 */ always @(posedge clk) if (1'b1) \data[18]  <= 1'b0 ? 1'b0 : n68;
/* FF  1 18  5 */ assign n24 = n69;
/* FF  1 27  4 */ assign n46 = n70;
/* FF  1 14  6 */ assign n16 = n71;
/* FF  1 21  4 */ assign n32 = n72;
/* FF  1 24  2 */ assign n41 = n73;
/* FF  1 21  3 */ assign n31 = n74;
/* FF  1 30  1 */ assign n51 = n75;
/* FF  1 22  3 */ assign n35 = n76;
/* FF  1 22  7 */ assign n36 = n77;
/* FF  1 16  1 */ assign n19 = n78;

endmodule

